settings.title = inställningar