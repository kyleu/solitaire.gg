general.number.one = ett
general.number.two = två
general.number.three = tre
general.number.four = fyra
general.number.five = fem
general.number.six = sex
general.number.seven = sju
general.number.eight = åtta
general.number.nine = nio
general.number.ten = tio
general.number.eleven = elva
general.number.twelve = tolv
options.resume = Återupptag spelet
options.resign = Avgå
options.redeal = Ny affär
options.same.deal = Samma Deal
options.winnable = Winnable Deal
settings.title = inställningar
settings.disclaimer = Jag jobbar på inställningssidan.
help.title = {0} Hjälp
help.about = Detta är {0}.
help.privacy.policy = {0} Sekretesspolicy
help.general = Hjälp för {0}.
help.play.now = Spela nu
help.also.known.as = Också känd som
help.objective = Mål
help.deck = Däck
help.layout = Layout
help.original.game = Original Spel
help.related.games = Relaterade spel
help.web.resources = Webresurser
help.rank.match.rule.none = ingen
help.rank.match.rule.up = en rang högre
help.rank.match.rule.down = en rang lägre
help.rank.match.rule.equal = samma rang
help.rank.match.rule.up.or.down = en rang lägre eller högre
help.rank.match.rule.up.by.2 = två nivåer högre
help.rank.match.rule.down.by.2 = två nivåer lägre
help.rank.match.rule.up.by.3 = tre nivåer högre
help.rank.match.rule.down.by.3 = tre rader lägre
help.rank.match.rule.up.by.4 = fyra nivåer högre
help.rank.match.rule.down.by.4 = fyra nivåer lägre
help.rank.match.rule.up.by.pile.index = en rang högre för den första högen, två högre för den andra och så vidare,
help.rank.match.rule.any = någon rang
help.suit.match.rule.none = ingen
help.suit.match.rule.same.suit = samma kostym
help.suit.match.rule.different.suit = en annan kostym
help.suit.match.rule.same.color = samma färg
help.suit.match.rule.alternating.color = en annan färg
help.suit.match.rule.any = någon kostym
help.fill.empty.with.any = En tom hög kan fyllas med vilket kort som helst.
help.fill.empty.with.none = En tom hög kan inte fyllas.
help.fill.empty.with.rank = En tom hög kan fyllas med någon {0}.
help.fill.empty.with.rank.until.stock.empty = En tom hög kan fyllas med någon {0} tills lagret är tomt.
help.fill.empty.with.high.rank.or.low.rank = En tom hög kan fyllas med någon {0} eller {1}.
help.fill.empty.with.sevens = En tom hög kan fyllas med några sju.
help.victory.condition.all.but.four.on.foundation = Placera alla utom fyra kort på stiftelsen.
help.victory.condition.all.on.foundation = Placera alla kort på fundamentet i följd.
help.victory.condition.all.on.foundation.or.stock = Placera alla kort på fundamentet eller lagret.
help.victory.condition.all.on.tableau.sorted = Sortera alla kort på bordet så att var och en är {0} och {1}, eller flytta dem till grunden.
help.victory.condition.none.in.pyramid = Ta bort alla kort från pyramiden.
help.victory.condition.none.in.stock = Ta bort alla kort från lagret och avfallet.
help.victory.condition.pairs.sr = Ta bort alla par med lika stora rader.
help.victory.condition.pairs.srsc = Ta bort alla par med samma räcker och samma färg.
help.victory.condition.pairs.ss = Ta bort alla par med samma kostym.
help.victory.condition.pairs.9-or-10jqk = Ta bort alla par som lägger till nio och alla Nines, Tens, Jacks, Queens och Kings.
help.victory.condition.pairs.10-or-10JQK-pairs = Ta bort alla par som lägger till tio, par Jacks, Queens par och Kings par.
help.victory.condition.pairs.10-or-10JQK = Ta bort alla par som lägger till tio, och alla Tens, Jacks, Queens och Kings.
help.victory.condition.pairs.10-or-four-10JQK = Ta bort alla par som lägger till tio, och alla uppsättningar av Tio, Jacks Queen och King.
help.victory.condition.pairs.11-or-JQK-pairs = Ta bort alla par som lägger till elva och alla par av Jacks, Queens, and Kings.
help.victory.condition.pairs.11-or-Jpair-or-QK = Ta bort alla par som lägger till elva, alla par av Jacks, och alla Queen / King-par.
help.victory.condition.pairs.11-or-JQK = Ta bort alla par som lägger till elva och alla Jacks, Queens och Kings.
help.victory.condition.pairs.ss-11-or-JQK = Ta bort alla samma kostympar som lägger till elva, och alla Jacks, Queens och Kings.
help.victory.condition.pairs.12-or-QK = Ta bort alla par som lägger till tolv, och alla Queens och Kings.
help.victory.condition.pairs.13-or-K = Ta bort alla par som lägger till 13 och alla Kings.
help.victory.condition.pairs.14 = Ta bort alla par som lägger till 14.
help.victory.condition.pairs.15-or-10JQK = Ta bort alla par som lägger till 15, och alla uppsättningar av Tio / Jack / Queen / King.
help.victory.condition.pairs.15-or-A-pair = Ta bort alla par som lägger till 15 och alla esspar.
help.victory.condition.pairs.15-or-four-10JQK = Ta bort uppsättningar som lägger till femton, och uppsättningar av alla fyra Tens, Jacks, Queens och Kings.
help.victory.condition.pairs.17-or-A23 = Ta bort alla par som lägger till 17, och alla uppsättningar av Ace / Two / Three.
help.victory.condition.pairs.face-and-three-that-add-to-18 = Ta bort alla uppsättningar av ett ansikte kort och tre andra som lägger till 18.
help.victory.condition.pairs.cr = Ta bort alla par med varandra följande rader.
help.victory.condition.pairs.cr-or-AK = Ta bort alla par med varandra i rad eller Ace / King.
help.victory.condition.pairs.cr-or-sr = Ta bort alla par med varandra i följd eller lika med varandra.
help.deck.single.standard = Ett standarddäck med {0} kort.
help.deck.single.oddranks = Ett däck med {0} kort med ledningar {1}.
help.deck.single.oddsuits = Ett däck med {0} kort med passar {1}.
help.deck.single.oddranksandsuits = Ett däck med {0} kort med hjälp av röster {1} och kostymer {2}.
help.deck.multiple.standard = {0} standarddäck totalt {1} kort.
help.deck.multiple.oddranks = {0} täcker totalt {1} kort med hjälp av ledningar {2}.
help.deck.multiple.oddsuits = {0} täcker totalt {1} kort med kostymer {2}.
help.deck.multiple.oddranksandsuits = {0} täcker totalt {1} kort med hjälp av röster {2} och kostymer {3}.
help.piles.single = En enda {0} hög.
help.piles.single.cards.empty = En enda tom {0} hög.
help.piles.single.cards.single = En enda {0} hög med ett initialkort.
help.piles.single.cards.multiple = En enda {0} hög med {1} initialkort.
help.piles.multiple = {0} {1} högar.
help.piles.multiple.cards.empty = {0} tomma {1} högar.
help.piles.multiple.cards.single = {0} {1} högar med ett initialkort som delas ut till dem.
help.piles.multiple.cards.single.each = {0} {1} högar med ett initialkort behandlat till vardera.
help.piles.multiple.cards.multiple = {0} {1} högar med {2} initialkort behandlade till dem.
help.piles.multiple.cards.multiple.each = {0} {1} högar med {2} initialkort behandlade till vardera.
help.piles.multiple.cards.pile.index = {0} {1} högar med ett kort som delas till första stapeln, två till andra, och så vidare.
help.piles.multiple.cards.rest.of.deck = {0} {1} högar med resten av korten i däcket som behandlas dem.
help.piles.multiple.cards.custom = {0} {1} högar med ett anpassat antal kort som delas ut till dem.
help.stock.cards.shown = {0} kort är synliga.
help.stock.cards.dealt.single = ett kort
help.stock.cards.dealt.multiple = {0} kort
help.stock.cards.dealt.fewer.each.time = tre kort, då färre varje gång,
help.stock.deal.to.foundation = När den väljs, handlar {0} till varje grundhög.
help.stock.deal.to.manually = Flytta manuellt kort från lageret.
help.stock.deal.to.never = Inga kort kan flyttas.
help.stock.deal.to.reserve = När det väljs, handlar {0} till varje reservpinne.
help.stock.deal.to.tableau = När den väljs, handlar {0} till varje tabellauhög.
help.stock.deal.to.tableau.first.set = När den väljs, handlar {0} till varje tabellau hög i den första uppsättningen.
help.stock.deal.to.tableau.if.none.empty = När det väljs, handlar {0} till varje tabellau hög om inget är tomt.
help.stock.deal.to.tableau.empty = När den väljs, handlar {0} till varje tom tabellhög.
help.stock.deal.to.tableau.non.empty = När den väljs, handlar {0} till varje icke-tom tabellauhög.
help.stock.deal.to.waste = När det väljs, handlar {0} till avfallet.
help.stock.deal.to.waste.or.pair.manually = När den väljs, handlar {0} till avfallet, eller kopplas manuellt.
help.stock.max.deals.single = Endast ett enda pass genom lageret är tillåtet.
help.stock.max.deals.multiple = Upp till {0} passerar genom lagret.
help.stock.max.deals.unlimited = Beståndet har obegränsade förlossningar.
help.waste.playable.cards.all = Alla kort kan flyttas från {0}.
help.waste.playable.cards.top = Det övre kortet kan flyttas från {0}.
help.foundation.lowrank.any = Alla kort kan flyttas till någon tom {0} hög.
help.foundation.lowrank.ascending = En Ace kan spelas den första {0} högen, en två på den andra och så vidare.
help.foundation.lowrank.first.becomes.base = Det första kortet som spelas till {0} blir baskortet för andra.
help.foundation.lowrank.specific = Alla {1} kan spelas till någon tom {0} hög.
help.foundation.initial.restriction.specific.color.unique.suits = Varje stapel måste startas med ett {0} kort och vara en unik kostym.
help.foundation.initial.restriction.specific.suit = Varje stapel måste startas med ett {0} kort.
help.foundation.initial.restriction.unique.colors = Varje stapel måste startas med en unik färg.
help.foundation.initial.restriction.unique.suits = Varje stapel måste startas med en unik kostym.
help.foundation.build.none = Inga kort kan byggas på ett kort i en {0} hög.
help.foundation.build.rank.and.suit.match.rules = Ett kort kan byggas på ett kort i en {0} hög om det är {1} och {2}.
help.foundation.wrap.ranks = En {0} kan spelas på en {1}, fortsätter sekvensen.
help.foundation.cards.shown = {0} kort är synliga.
help.foundation.move.complete.sequences.only = Kompletta sorterade sekvenser av kort kan flyttas en tom {0} hög.
help.tableau.unique.ranks = Pålarna hanteras på ett sådant sätt att inga två kort i samma stapel har samma rang.
help.tableau.cards.face.down.all.but.one = Toppkortsen på varje hög är vänd uppifrån.
help.tableau.cards.face.down.none = Alla kort är vända uppåt.
help.tableau.cards.face.down.single = Allt utom det första kortet i varje hög är vänd uppifrån.
help.tableau.cards.face.down.multiple = Alla utom de första {0} korten i varje hög är vända uppåt.
help.tableau.cards.face.down.even.numbered = Varje udda numrerat kort vänds uppifrån.
help.tableau.cards.face.down.odd.numbered = Varje jämnt numrerat kort vänds uppåt.
help.tableau.build.none = Inga kort kan byggas på ett kort i en {0} hög.
help.tableau.build.rank.and.suit.match.rules = Ett kort kan byggas på ett kort i en {0} hög om det är {1} och {2}.
help.tableau.move.stacks.none = Inga kort kan flyttas från {0} högar.
help.tableau.move.stacks.rank.and.suit.match.rules = Stackar av kort kan flyttas från en {0} hög om de är {1} och {2}.
help.pyramid.rows.single = en enda rad
help.pyramid.rows.multiple = {0} rader
help.pyramid.type.standard = En standard {0} med {1} (den övre raden har bara ett kort, två i nästa och så vidare).
help.pyramid.type.inverted = En inverterad {0} med {1} (den nedre raden har bara ett kort, två i nästa och så vidare).
help.pyramid.wrap.ranks = En ess kan spelas på en kung, fortsätter sekvensen.
help.pyramid.build.none = Inga kort kan byggas på denna {0}.
help.pyramid.build.rank.and.suit.match.rules = Ett kort kan byggas på detta {0} om det är {1} och {2}.
help.pyramid.move.stacks.none = Inga kort kan flyttas från {0}.
help.pyramid.move.stacks.rank.and.suit.match.rules = Kort kan flyttas från detta {0} om de är {1} och {2}.
rules.aceofhearts.description = Alla kort måste byggas på en enda grundpelare i denna Thomas Warfield-uppfinning.
rules.acesandkings.description = Bygg upp på en grund, ner på den andra, men bygg inte alls på bordauen.
rules.aceyandkingsley.description = En variation av ^ acesandkings ^ som börjar med en ess eller en kung som behandlas till varje stiftelse.
rules.acme.description = En svår variant av ^ canfield ^ där du bygger i kostym, kan inte flytta sekvenser och bara få två passeringar genom lagret.
rules.acquaintance.description = En variation av ^ auldlangsyne ^ föreslog av Michael Keller som lägger till något intresse genom att tillåta två lösningar.
rules.adelaide.description = Denna tvådels-kabal gör det möjligt att flytta osorterade staplar, som i ^ yukon ^.
rules.agnesbernauer.description = En variation på ^ klondike ^ med sju reserver.
rules.agnessorel.description = En variation på ^ klondike ^ där kort behandlas direkt på bordet som i ^ spider ^.
rules.alaska.description = En något svårare variant av ^ yukon ^ där du kan bygga upp eller ner, men måste bygga i samma färg.
rules.alexanderthegreat.description = Thomas Warfields mer utmanande variation av ^ Cloverleaf ^.
rules.alexandria.description = En tre-däckversion av ^ tjuvesofegypt ^ uppfunnad av Thomas Warfield.
rules.algiers.description = En tredäcksvariant av ^ karthage ^.
rules.alibaba.description = En-däckvariation av ^ fyrtiondag ^ där du kan flytta sekvenser av kort ihop istället för bara en i taget.
rules.allinarow.description = En variation av ^ golf ^ utan ett lager.
rules.alternate.description = En variation av ^ sirtommy ^ där grunden är byggd i alternativ färg, halv uppåt, halv nedåt.
rules.alternations.description = En variation av ^ utbyte ^ som har samma 7 till 7 tabellau med alternativa kort med framsidan nedåt, men där du bygger in alternativa färger.
rules.alternative.description = Denna relativitet av ^ klöverbladet ^ tillåter inte att mellanslag fylls men tillåter en återlösning.
rules.americancanister.description = En svår variant av ^ canister ^ med byggnad av alternativa färger.
rules.americantoad.description = En enkel tvådäcksvariant av ^ canfield ^.
rules.antares.description = Thomas Warfields kombination av ^ freecell ^ och ^ scorpion ^ delar in tabellen i två halvor, en där vi bygger i alternativa färger och flyttar kort med FreeCell regler, en där vi bygger i samma kostym och flyttar med Scorpions regler.
rules.ants.description = Liksom fyra parallella ^ golf ^ -spel
rules.anubis.description = En variation av ^ doublepyramid ^ med tre avfallspiller.
rules.apophis.description = ^ pyramid ^ spelas med tre avfallspiller.
rules.applegate.description = Detta spel har likheter med både ^ spider ^ och ^ yukon ^ och kan vara en äldre version av ^ scorpion ^
rules.arabella.description = En tre-deck ^ spider ^ / ^ klondike ^ blandar sig med ^ ladyjane ^ av Thomas Warfield.
rules.arizona.description = En lättare variation av ^ wildflower ^ där du kan flytta sekvenser oavsett kostym.
rules.assembly.description = Kostymer spelar ingen roll alls i detta enkla lilla solitaire spel.
rules.astrocyte.description = Ett komprimerat spel av ^ spider ^ med fyra celler.
rules.athena.description = A ^ klondike ^ -variation med en rektangulär startbordsbana i vilken kort växlar uppifrån och nedåt.
rules.auldlangsyne.description = Ett gammalt solitaire spel där ingen byggnad är tillåten på bordet.
rules.auntmary.description = En svår ^ klondike ^ variant där bordet innehåller en mindre stapel men alla kort är vända uppåt.
rules.australian.description = En variation av ^ klondike ^ som tillåter att icke-toppkort flyttas (med korten ovanpå dem) som i ^ yukon ^.
rules.backbone.description = Ett svårt spel av viktorianskt ursprung med en gaffelreserv
rules.bakers.description = En föregångare till ^ freecell ^ uppfunnad av C. L. Baker.
rules.bakersdozen.description = Ordna om de tretton tableau-staplarna för att frigöra kort till grunden genom att flytta ett kort åt gången.
rules.bakerstwodeck.description = En två-däckversion av ^ bakare ^ -spel.
rules.balcony.description = Liknande ^ canfield ^, men grundarna är uppbyggda i alternativa färger kan reservkort endast spelas till grunden, och tomma utrymmen är autofyllda från lagret.
rules.barricadea.description = Ett enkelt spel där vi bygger oberoende av kostym på både bordau och foundation och som använder ett lager men inte ett slöseri.
rules.barricadeb.description = En lättare, men fortfarande mycket svår, modifiering av ^ block ^ uppfunnet av Richard Mechen och Thomas Warfield.
rules.bastion.description = ^ fästning ^ med celler.
rules.bath.description = A ^ freecell ^ variant där utrymmen endast kan fyllas av kungar och det finns bara två celler.
rules.batsford.description = Ett två-deck ^ klondike ^ spel med en speciell reserv som kan lagra upp till tre kungar.
rules.batsfordagain.description = En variation av ^ batsford ^ med en redeal.
rules.bavarian.description = Thomas Warfields enklare version av ^ tyska ^ tålamod med några extra tabellau kolumner.
rules.bearriver.description = A ^ fan ^ variation där du kan bygga upp och ner i kostym, men är begränsad till tre kort per hög.
rules.beehive.description = I detta ^ lagerhus ^ variant bygger och tar vi bort staplar av fyra kort med samma rang.
rules.beehivegallery.description = Det här är bara ^ beehive ^ med ett annat användargränssnitt: alla kort som normalt skulle startas i lagret blinkas uppåt med de som normalt skulle kunna spelas om du gick igenom lagret tre åt gången automatiskt
rules.beetle.description = En variant av ^ spider ^ där alla kort hanteras uppåt.
rules.beleagueredcastle.description = Ett utmanande spel med enkla regler.
rules.beleagueredfortress.description = En variation av ^ fästning ^ med en tolv-kort reserv, från vilken alla kort är spelbara.
rules.bigapple.description = En svår variant av ^ newyork ^ med tre celler i stället för tre avfallspiller, men där staplar kan flyttas.
rules.bigbertha.description = Denna tvådäcksversion av Kingalbert ^ som har 14 reservkort som är alla spelbara och en separat grundval som du kan lägga på alla kungarna.
rules.bigforty.description = En-däckvariant av ^ fyrtiofier ^ som tillåter stapelrörelser.
rules.bigfreecell.description = En rakt framåt två-däckversion av ^ freecell ^.
rules.bigharp.description = En två-däck ^ klondike ^ -variation som är annorlunda än ^ harp ^ på flera sätt, utan att verkligen vara så mycket större.
rules.bigspider.description = En tre-däckversion av ^ spider ^.
rules.binarystar.description = Thomas Warfields tvådäcksversion av ^ blackhole ^ har två grundpelare.
rules.bisley.description = Ett spel att bygga upp och ner på bordet.
rules.blackhole.description = Liksom ^ allinarow ^, detta är en variation av ^ golf ^ utan ett lager.
rules.blackwidow.description = En lättare variant av ^ spider ^ där du får flytta sekvenser även om de inte är alla ena kostym.
rules.blindalleys.description = A ^ klondike ^ variant med en fyrkantig tabellau, som skiljer sig från ^ passeul ^ endast i antalet passerar genom det tillåtna däcket.
rules.block.description = Ett nästan oväldigt svårt två-däck spel som får sitt namn från det faktum att det rutinmässigt blockerar.
rules.blockade.description = Ett enkelt spel som börjar långsamt och slutar med en blomstring.
rules.blockten.description = Ett spel av ren tur där du kan ta bort par som lägger till tio, eller par av ansikte kort, men inte tiotals.
rules.blondesandbrunettes.description = En variant av ^ signora ^ där grundbaskortet bestäms av ett kort som delas in.
rules.bobby.description = En variation av ^ robert ^ med en andra foundation stapel för att underlätta, men inte mycket lättare.
rules.boulevard.description = Ingen byggnad på bordet, tre reservpeler och stiftelser som byggs upp genom två.
rules.boxfan.description = A ^ fan ^ variant med byggnad med alternativ färg.
rules.boxkite.description = Tableaus byggs upp eller ner, halva grundarna byggs upp, halva bygga ner.
rules.brazilian.description = I denna två-däck ^ klondike ^ -varianten från Brasilien handlar du om bordläggningen istället för att ha en avfallspole.
rules.breakwater.description = En lättare variant av ^ utbyte ^, där vi bygger oberoende av kostym.
rules.brigade.description = En lättare variation av ^ flowergarden ^ med fler bordau högar med färre kort och ess som börjar på grunden.
rules.brisbane.description = Precis som ^ yukon ^, men startlayouten är lite annorlunda och du bygger oberoende av kostym.
rules.bristol.description = Ett spel med tre spillpiller uppfunna av Albert Morehead och Geoffrey Mott-Smith.
rules.britishcanister.description = En svår version av ^ canister ^ som går tillbaka till 1890-talet.
rules.brownrecluse.description = Denna ^ spindel ^ variant av Thomas Warfield har ett lager och en avfallspål.
rules.bucket.description = A ^ canister ^ -variation som slutar ser ganska som ^ freecell ^ utan cellerna.
rules.buffalobill.description = I denna lätta variant av ^ littlebillie ^, av David Parlett, finns det fler fans och reservcellerna börjar tomma, men det finns inga lösningar.
rules.bunker.description = Bygg upp oavsett kostym för att försöka få alla kort på bordet.
rules.bureau.description = Detta spel har regler som liknar ^ klondike ^, förutom att du bygger grunden i alternativa färger och inte kan fylla utrymmen i tabellau.
rules.busyaces.description = Ett ganska enkelt spel som går tillbaka till 1939. Tolv bordaustackar med ett kort betyder att du enkelt kan få massor av tomma utrymmen att arbeta med.
rules.calculation.description = I grunden liknar ^ sirtommy ^, men mycket mer komplext att spela eftersom varje fundament staplar framåt med ett annat steg.
rules.canfield.description = Ett gammalt kasinospel där huset vanligtvis vinner.
rules.canfieldgallery.description = Det här är bara ^ canfield ^ med ett annat användargränssnitt: Alla kort som normalt skulle startas i aktien blinkas uppåt med de som normalt skulle kunna spelas om du gick igenom lagret tre åt gången automatiskt
rules.canfieldrush.description = A ^ canfield ^ variant där kort behandlas av tre i första passet, två gånger i andra och en-i-ett-tiden i det sista.
rules.canister.description = Ännu ett generiskt solitaire spel, med alla kort handlade fram och inga lager.
rules.caprice.description = Bygg upp eller ner i kostym och lagerhandlar till bordau.
rules.captivequeens.description = En enkel och hjärnlös variation av ^ sixesandsevens ^ också känd som \
rules.carlton.description = En svår två-däck ^ klondike ^ -variation.
rules.carousel.description = Ett tvådäcksspel med separata fundament för ess, evens och odds.
rules.carpet.description = En lätt match med tjugo reservposter och ingen byggnad.
rules.carthage.description = En två-däck spel där du hanterar reserverna och bygger på bordet.
rules.cassim.description = En version av ^ alibaba ^ med en mindre tabellau och en oändlighet av förlossningar.
rules.castile.description = En öppen variant av ^ bristol ^ uppfunnad av Thomas Warfield.
rules.castlemount.description = En tre-däckversion av ^ beleagueredcastle ^ uppfunnet av Thomas Warfield.
rules.castleofindolence.description = Thomas Warfields anpassning av ett 19th century-spel som först beskrivs i George A. Bonaventures 1932-bok med solitaire-spel.
rules.castlesend.description = En något annorlunda version av ^ schackbräda ^ med en kort med två kort.
rules.castlesinspain.description = En variant av ^ bakersdozen ^ som gör det möjligt att fylla i mellanslag med något kort och där vi bygger in alternativa färger.
rules.castoutnines.description = En svår variant av ^ deuces ^ eller ^ busyaces ^ där inga kort redan finns på grunden och det finns bara sju tableau-staplar.
rules.ceilingfan.description = En lättare variant av ^ fan ^ där du bygger in alternativa färger.
rules.celleleven.description = En tre-däckversion av ^ freecell ^.
rules.challengefreecell.description = En version av ^ freecell ^ uppfunnad av Thomas Warfield där ess och twos alltid ligger på botten av de åtta staplarna.
rules.chameleon.description = Om ^ canfield ^ inte var tillräckligt svårt för dig, är det här en version med bara tre bordsskenor.
rules.chateau.description = En två-deck ^ beleagueredcastle ^ variant.
rules.chelicera.description = En variation på ^ scorpion ^ uppfunnad av Erik den Hollander, där vi fyller utrymmen med tre kort från lageret istället för att hantera lageret.
rules.cheops.description = En variant av ^ pyramiden ^ där du tar bort par av kort med lika eller i följd rader
rules.chequers.description = Det här spelet har tjugofem tableau högar där du kan bygga upp eller ner, och du bygger upp på hälften av fundamenten och ner på de andra.
rules.chessboard.description = En mer intressant variation av ^ fästning ^ där du väljer baskortet.
rules.chinaman.description = A ^ klondike ^ variant där vi bygger olika drag.
rules.chinese.description = Denna ^ skorpion ^ -variation har en annan layout, ett mindre lager och låter kort flyttas till stiftelsen en åt gången.
rules.chinesefreecell.description = En version av ^ freecell ^ spelas med endast tre drag.
rules.chineseklondike.description = En tre-färgversion av ^ klondike ^.
rules.chinesespider.description = En tre-kostymversion av ^ spider ^.
rules.cicely.description = En variation av ^ turnering ^ och ^ kingsdowneights ^ där du kan bygga upp och ner på bordet.
rules.circleeight.description = Flytta alla kort till bordet för att vinna detta spel, men du kan inte flytta ett kort när det är på bordet.
rules.citadel.description = En lättare variation av ^ beleagueredcastle ^ där kort flyttas till stiftelsen under affären.
rules.cleopatra.description = Thomas Warfields variant av ^ fortythieves ^ med en pyramidformad tableau.
rules.cloverleaf.description = En lätt spel uppfunnad av Thomas Warfield där du bygger upp eller ner på bordet, bygger två grundpelare upp och två bygger ner.
rules.colonel.description = En variation av ^ signora ^ uppfunnit av Thomas Warfield där vi byggde i samma kostym istället för växlande färger.
rules.colorado.description = Ett spel där kort kan staplas godtyckligt på 20 bordålar.
rules.congress.description = Detta har likheter med ^ fyrtiondag ^, men utrymmen i bordet får endast fyllas av avfallet.
rules.contradance.description = En variation av ^ sixesandsevens ^ som är lika hjärnlös som ^ captivequeens ^, men kräver mycket större lycka att någonsin vinna.
rules.cornelius.description = En version av ^ fyrtiondag ^ som tillåter att icke-bästa kort spelas (flytta vilka kort som är ovanpå dem tillsammans med dem) som i ^ yukon ^.
rules.corners.description = Denna helt tanklösa variant på ^ czarina ^ tillåter ingen byggnad på bordau men tillåter tre passerar genom beståndet.
rules.cornersuite.description = Det här ganska lätta spelet liknar en däckversion av ^ kongress ^, förutom att tabellen börjar tom.
rules.corona.description = Ett spel som liknar ^ fyrtiondag ^ där utrymmen är autofyllda från avfall och lager.
rules.countess.description = A ^ canfield ^ -variation med fyra reserver.
rules.courtyard.description = En variation av ^ upptagssatser ^ som ökar svårigheten genom att autofyllning av tomma bordutrymmen avfall och lager.
rules.coyote.description = En något lättare, men fortfarande svår, variation av ^ acme ^ i vilken sekvenser kan flyttas.
rules.crescent.description = Ett dubbelriktat byggnadsspel där du kan rotera kort i staplarna tre gånger.
rules.crescentfour.description = En lättare variation av ^ crescent ^ som tillåter en extra rotation.
rules.crisscross.description = En variation av ^ simplepairs ^ som kräver en mycket stor dos av ren tur att vinna.
rules.cromwell.description = Ett tvådäcksspel med 26 tableau högar och en rita.
rules.cruel.description = Ett spel där du kan redovisa tabellen så ofta du vill, så länge du kan ta bort minst ett kort mellan erbjudanden.
rules.czarina.description = En variation på ^ fourseasons ^ där utrymmen fylls automatiskt från beståndet.
rules.darkpyramid.description = En version av ^ pyramiden ^ där korten behandlas nedåt.
rules.darwin.description = En tre-däckversion av ^ australian ^ Solitaire, som är ett kors mellan ^ yukon ^ och ^ klondike ^.
rules.demon.description = En två-däckversion av ^ canfield ^, inte lika lätt som ^ doublecanfield ^.
rules.demonfan.description = En väldigt lätt spel där du bygger ner i alternativa färger och får sex redovisningar.
rules.demonsandthieves.description = I det här spelet är uppdelningen uppdelad i två halvor, en halv där du spelar med ^ canfield ^ -regler och en halv där du spelar med ^ fyrtiofire regler.
rules.deuces.description = En svårare variant av ^ uppspelning ^ med färre bordauhögar.
rules.deucesandqueens.description = En variation på ^ acesandkings ^ där byggnaden är tillåten på bordet.
rules.diavolo.description = A ^ klondike ^ variant med fyra grundstaplar som byggs ett kort åt gången, medan de andra fyra behöver slutförda sekvenser.
rules.dieppe.description = En variation på ^ kongressen ^ där staplar kan flyttas, kan blanketter fyllas med vilket kort som helst och tre rader kort behandlas initialt.
rules.dimes.description = En variation på ^ deuces ^ med färre tableau högar.
rules.diplomat.description = En variation på ^ kongress ^ eller ^ fyrtiondag ^.
rules.dnieper.description = Exakt som ^ kiev ^ men lite lättare eftersom kungar kan spelas på ess.
rules.dorothy.description = En annan hjärnlös variation av ^ captivequeens ^ och ^ sixesandsevens ^ med separata fundament för odds, evens och face cards.
rules.doubleacesandkings.description = En fyrdäcksversion av ^ acesandkings ^ uppfunnad av Thomas Warfield.
rules.doublecanfield.description = En två-däckversion av ^ canfield ^, mycket mycket lättare än det ursprungliga spelet.
rules.doubledot.description = En lätt spel där du bygger upp två på grunden, och ner vid två på bordet.
rules.doubleeasthaven.description = En tvådäcksversion av ^ easthaven ^.
rules.doublefourteens.description = En två-däckversion av ^ fourteenout ^.
rules.doublefreecell.description = Thomas Warfields tvådäcksversion av ^ freecell ^.
rules.doublegoldrush.description = En tvådäcksversion av ^ goldrush ^.
rules.doublejane.description = En fyra däck ^ spider ^ / ^ klondike ^, liknande ^ ladyjane ^.
rules.doubleklondike.description = En två-däckversion av ^ klondike ^.
rules.doublelimited.description = En fyrdäcksversion av ^ begränsad ^.
rules.doubleminerva.description = Thomas Warfields tvådäcksversion av ^ minerva ^.
rules.doublepyramid.description = Thomas Warfields tvådäcksversion av ^ pyramiden ^.
rules.doublerail.description = A ^ fortythieves ^ variation där vi bygger oberoende av kostym och kan flytta staplar.
rules.doublerussian.description = En två-däckversion av ^ russian ^ solitaire.
rules.doublescorpion.description = En enkel tvådäcksvariant av ^ scorpion ^ där alla kort redan behandlas i början.
rules.doubleseatowers.description = En tvådäcksversion av ^ freecell ^ -varianten känd som ^ sitsar ^.
rules.doublesignora.description = En fyrdäcksversion av ^ signora ^ uppfunnad av Thomas Warfield.
rules.doublestorehouse.description = En tvådäcksversion av ^ lagerhus ^.
rules.doubletcell.description = En kombination mellan ^ dubblets ^ och ^ freecell ^.
rules.doubletrigon.description = En två-deck version av ^ trigon ^ eller kanske en version av ^ doubleklondike ^ med byggnad i kostym.
rules.doublets.description = Ett liknande spel till ^ simplepairs ^.
rules.doubleyukon.description = En tvådelsvariation av ^ yukon ^
rules.dover.description = Denna tvådäcksversion av ^ bristol ^ har fortfarande tre avfallspeler, men grundpinnar måste byggas upp i kostym och tomma bordutrymmen kan fyllas, men endast från avfallet.
rules.dragon.description = En variation av ^ kinesiska ^ där du bygger i samma kostym.
rules.easthaven.description = En en-däck korsning mellan ^ spider ^ och ^ klondike ^.
rules.eclipse.description = En variant av ^ waningmoon ^, där sekvensen rör sig är tillåtet och kort behandlas till bordau istället för till en avfallspole.
rules.eightbyeight.description = Bygg oavsett kostym på en 8x8 bordau för att få dina kort på de åtta grundarna.
rules.eighteens.description = Ett spel där du tar bort singleton ess, eller uppsättningar som består av ett ansikte kort med tre andra kort som lägger till arton.
rules.eightoff.description = A ^ freecell ^ variation med fler celler, men där du bara kan bygga ner i samma färg
rules.eighton.description = En hårdare variation av ^ eightoff ^ där esserna börjar på bottnen av pålarna.
rules.eightsdown.description = A ^ busyaces ^ variant uppfunnad av Thomas Warfield, där grunden bygger ner från åtta.
rules.eightythieves.description = En mycket svår fyrdäcksversion av ^ fortythieves ^ av Thomas Warfield.
rules.elba.description = En variant av fyrtiofem med ^ klondike ^ -liknande byggregler.
rules.elevens.description = En uppsättning avlägsnande uppsättningar av kort som lägger till 15 eller uppsättningar som innehåller tio genom kungen.
rules.eleventriangle.description = En något enklare version av ^ triangle ^ där vi tar bort par som lägger till elva.
rules.eliminator.description = Ett enkelt ^ golf ^ -liknande spel med sex stiftelser.
rules.emperor.description = En svårare version av ^ rankandfile ^ där endast enskilda kort kan flyttas ..
rules.empressofitaly.description = En fyrdäcksversion av ^ blondesandbrunettes ^ uppfunnad av Thomas Warfield.
rules.endlessharp.description = En variation av Big Harp som tillåter obegränsad förlossning.
rules.ephemeralfreecell.description = Ephemeral FreeCell är som standard ^ freecell ^, förutom att en av cellerna kommer att försvinna efter det första användningen.
rules.escalator.description = Dekonstruera en pyramid genom att bygga upp eller ner på en enstaka stapel.
rules.eternaltriangle.description = En ganska svår två-däck ^ klondike ^ -variation.
rules.evenandodd.description = En-däckversion av ^ boulevard ^.
rules.exiledkings.description = En svårare variation av ^ citadel ^ där utrymmen endast kan fyllas av kungar.
rules.fairmaids.description = En variation av ^ willothewisp ^ där vi bygger in alternativa färger.
rules.fallingstar.description = En svåra ^ signora ^ -variation med en mindre tabellau-stapel och en förutbestämd grundbas.
rules.famousfifty.description = En svår ^ förtythieves ^ -variation som börjar med ett extra kort på varje bordauhög.
rules.fan.description = Det ursprungliga Fan-spelet innebär att bygga i klädsel på arton tableau-staplar.
rules.farmerswife.description = En variation av ^ treblindmus ^ där vi bygger in alternativa färger som i ^ scorpiontail ^.
rules.father.description = Denna variation av ^ farfar ^ av Thomas Warfield lägger till svårigheter genom att minska antalet bordauhögar och lägger till strategi genom att eliminera automatisk fyllning av tomma utrymmen, men det är fortfarande ett ganska enkelt spel.
rules.fifteen.description = Bygg upp på en grund, nere på den andra.
rules.fifteenrush.description = Layouten är som ^ klondike ^, men du tar bort par som lägger till femton eller par esser.
rules.fifteens.description = Ett enkelt spel där du tar bort uppsättningar som lägger till 15 eller uppsättningar av fyra tiotals, fyra jacks, fyra drottningar eller fyra kungar.
rules.floradora.description = En två-däck variant av ^ thirtysix ^ med en extra fundament stapel för kungar, men ingen stack rör sig.
rules.flow.description = En lättare variation av ^ wavemotion ^ som tillåter att bygga på reserven.
rules.flowergarden.description = De sex staplarna av sex kort i bordau kallas \
rules.fly.description = En variation av ^ groda ^ där esserna börjar på grunden.
rules.forecell.description = En svensk föregångare till ^ freecell ^, ursprungligen en av många spel som heter \
rules.fortress.description = En klassisk och vanligtvis obestridlig förfader till ^ beleagueredcastle ^ där du kan bygga både upp och ner i bordet.
rules.fortressofmercy.description = En variant av ^ fästning ^ som låter dig få en \
rules.fortunesfavor.description = En extremt enkel, en-däckversion av ^ busyaces ^.
rules.fortyandeight.description = Två däck, fyrtio kort i bordet, åtta grundpinnar, bygga i samma kostym.
rules.fortybandits.description = En lättare variant av ^ fortythieves ^ där sekvenser kan flyttas.
rules.fortydevils.description = Thomas Warfields svåra kors mellan ^ rougeforty ^ och ^ ladycadogan ^.
rules.fortynine.description = Denna förtyndring ^ -variationen har nittio nio kort i en sju av sju tabellau.
rules.fortythieves.description = Liknande ^ fyrtiondag ^, men tableauen har fyrtio kort i tio staplar av fyra, och vi tillåter bara en att passera genom däcken.
rules.fortythieves3.description = En tre däckversion av ^ fortythieves ^ med en 12 av 4 bordau.
rules.fortythieves4.description = En fyra däckversion av ^ fortythieves ^ med en 14 av 6 bordau.
rules.fourbyten.description = A ^ freecell ^ -variation med massor av celler och inte så många tableau-staplar.
rules.fourleafclovers.description = En enstaka stapel är byggd oavsett kostym från ess till kung och sedan från ess till kung igen med hjälp av en bordau där du kan bygga både upp och ner.
rules.fourseasons.description = Ett enkelt lycko och färdighet där du flyttar kort en åt gången, staplar oavsett kostym.
rules.foursup.description = Thomas Warfield skapade detta spel som en fortsättning på serien som börjar med de traditionella spelen ^ busyaces ^ och ^ deuces ^.
rules.fourteenout.description = Ett intressant spel där du tar bort par som lägger till fjorton.
rules.fredsspider.description = I denna lätta variant på ^ spider ^, designad av Fred Lunde i Livonia, Michigan, behandlas kort upp och kan flyttas till stiftelsen ensam.
rules.freecell.description = Inventad av Paul Alfille, känd av Microsoft, erbjuder detta spel fyra tillfälliga lagringsceller som kan användas för att flytta kort.
rules.freecellduplex.description = En enkel tvådäcksversion av ^ freecell ^.
rules.freecellfourdeck.description = En fyrdäcksversion av ^ freecell ^ för dem som gillar att tillbringa lång tid att lösa en enda affär.
rules.freecellthreedeck.description = Ännu en tre-däckversion av ^ freecell ^.
rules.freefan.description = En enkel variant av ^ fan ^ med celler.
rules.friday.description = Ett paravlägsningsspel med en tvådelig tabellau, varav endast en är autofylld från lagret.
rules.frog.description = En relation av ^ sirtommy ^ med en reserv.
rules.gargantua.description = En två-däckversion av ^ klondike ^ uppfunnad av Albert Morehead och Geoffrey Mott-Smith.
rules.gaygordons.description = Ett par borttagning spel där du tar bort par som lägger till 11, Kings med Queens eller Jacks tillsammans.
rules.german.description = Ett konstigt och svårt spel där du måste bygga sekvenser på bordet, oavsett kostym.
rules.giant.description = A ^ missmilligan ^ variant utan en ficka men i vilken kort som helst kan spelas till ett tomt utrymme.
rules.gilbert.description = En udda ^ klondike ^ -variation med en uppsättning av fundament som bygger upp och en uppsättning byggnad.
rules.giza.description = Michael Kellers variant av ^ pyramiden ^ har en tabellau av kort istället för ett lager, vilket gör det till ett helt öppet spel.
rules.gloucestershire.description = En tvådäcksvariant av ^ flowergarden ^.
rules.goldmine.description = A ^ klondike ^ variation som börjar med en tom tabellau.
rules.goldrush.description = A ^ klondike ^ variation där antalet kort som behandlas till avfallet minskar med varje passering genom lagret.
rules.golf.description = Bygg upp eller ner på den enda stiftelsen för att ta kort av bordau, där ingen byggnad är tillåten.
rules.golfrush.description = En variant av ^ golf ^ spelade på med en ^ klondike ^ -stils tabellau.
rules.goodmeasure.description = En mycket svårare variation av ^ bakersdozen ^ med färre bordsfält.
rules.gotham.description = En lättare variant av ^ newyork ^ där vi bygger oberoende av kostym och samma kostym kan flyttas.
rules.grandfather.description = Ett spel med tjugo bordshögar, som alla kan hålla två kort.
rules.greattriangle.description = En svår tre-deck ^ klondike ^ -version av Thomas Warfield.
rules.groundsfordivorce.description = A ^ spider ^ -spel där kort inte behandlas för att tömma kolumner.
rules.gypsy.description = Ett kors mellan ^ spider ^ och ^ klondike ^.
rules.halfcell.description = ^ freecell ^ med endast två grundstaplar.
rules.harp.description = En två-däck ^ klondike ^ -variation.
rules.haystack.description = En svårare version av ^ nål ^ där endast 8 kort kan lagras i reserven.
rules.howtheyrun.description = En variation av ^ threeblindmice ^ uppfunnad av Erik den Hollander med två celler som ersätter tvåkortsreserven.
rules.hugespider.description = En fyrdäcksversion av ^ spider ^.
rules.hypotenuse.description = En version av ^ eternaltriangle ^ med några kort vänd nedåt.
rules.imperialguards.description = En version av ^ missmilligan ^ där tomma tabellutrymmen kan fyllas med något kort istället för kungar.
rules.incompatibility.description = A ^ spider ^ -spel där kort kan flyttas till grunden en åt gången och där kort inte behandlas för att tömma kolumner.
rules.indefatigable.description = Denna variation av ^ royalfamily ^ är i grunden densamma, men grunden bygger upp från ess och det görs ännu lättare med en extra redaktion.
rules.indian.description = En lätt match som liknar ^ förtytieven ^, förutom att det första kortet i varje stapel av 10 bordet 3 är vänd nedåt och kort kan spelas på någon annan kost än sin egen.
rules.inquisitor.description = Denna ^ ladyjane ^ -variation av Thomas Warfield kräver att du bygger i kostym, men ger dig en extra redovisning.
rules.insaneklondike.description = En variation av ^ klondike ^ med 32 däck.
rules.intelligence.description = En två-däckversion av ^ labellelucie ^.
rules.interchange.description = En extremt svår ^ förtythieves ^ variant med alternativa kort behandlades med ansiktet nedåt.
rules.invertedfreecell.description = Precis som ^ freecell ^ men vi limber upp våra hjärnor genom att bygga allt i motsatt riktning.
rules.irmgard.description = En variant av ^ gypsy ^ där du har en extra tabellau hög, men du kan bara fylla utrymmen med kungar.
rules.isabel.description = Ta bort kortpar av samma rang från en 13x4 bordläggning.
rules.jacksinthebox.description = En variation på ^ deuces ^ som har färre tableau högar men lägger till några celler.
rules.josephine.description = Liknande ^ fyrtiofier ^, förutom att du kan flytta sekvenser.
rules.jumboklondike.description = ^ klondike ^ spelas med en sex-kostym däck.
rules.junction.description = En variation av ^ singlerail ^ eller ^ doublerail ^ för fyra piquet decks.
rules.juvenile.description = Ett tvådäcksspel där du tar bort par som lägger till fjorton.
rules.kansas.description = Liksom ^ regnbåge ^ det här är en ^ canfield ^ -variant där du bygger oberoende av kostym, men det här är lite svårare eftersom du bara har tre bordbunkar.
rules.kiev.description = En version av ^ ukrainska ^ Solitaire där det finns ett lager av kort behandlade till en rektangulär bordau, vilket gör hela saken snarare ^ spider ^ ish.
rules.kingalbert.description = Detta spel, ett av flera spel, även känt som \
rules.kingcell.description = En variation av ^ freecell ^ där vi bygger ner oavsett kostym istället för av alternativ färg, och endast kungar kan spelas för att tömma tabellutrymmen
rules.kingdom.description = Ett spel där ingen byggnad är tillåten i bordet och kostymer ignoreras när man bygger upp bordau.
rules.kingsdowneights.description = Denna variation av ^ -turneringen ^ har en tabellau där du kan bygga av alternativ färg i stället för celler.
rules.kingsley.description = Reverse ^ klondike ^ som i teorin är inte svårare, men som visar sig svårt att linda huvudet om du är van vid att spela den omvänden.
rules.kingtut.description = En pyramidvariation där vi hanterar tre kort på en gång och har obegränsade förlossningar.
rules.klondike.description = Världens mest kända solitaire spel har en triangulär bordau där du bygger ner i växlande färger.
rules.klondikegallery.description = Världens mest kända solitaire spel spelade i galleri läge så alla lager kort är alltid synliga och de spelbara de är upptagna
rules.klondike1card.description = Världens mest kända solitaire spel har en triangulär bordau där du bygger ner i växlande färger.
rules.klondiketerritory.description = Ett kors mellan ^ flowergarden ^ och ^ klondike ^, något svårare än det liknande nordvästra territoriet spelet.
rules.knottynines.description = En svårare variant av trustytwelve ^.
rules.labellelucie.description = En klassisk solitaire där du bygger ner i kostym på bordet och kan redisera två gånger.
rules.ladybetty.description = Denna kusin av ^ sirtommy ^ kräver att du bygger stiftelsen i kostym, men ger dig två extra bordsskivor att arbeta med.
rules.ladycadogan.description = Thomas Warfields ^ rougeetnoir ^ variant där vi bygger oavsett kostym istället för i alternerande färger.
rules.ladyjane.description = En lätt två-deck ^ spider ^ / ^ klondike ^ blandning av Thomas Warfield.
rules.ladypalk.description = Liknande ^ diplomat ^, men tillåter att staplar flyttas och utrymmen kan bara fyllas av kungar.
rules.lafayette.description = A ^ canfield ^ variant med en grundbyggnad och en byggnad.
rules.lanes.description = En sex-av-tre-tabell spelade mycket som ^ klondike ^, men du kan inte flytta staplar.
rules.lasker.description = En version av ^ schackbräda ^ där sekvenser kan flyttas.
rules.leapyear.description = En fyra-däckversion av ^ auldlangsyne ^.
rules.lily.description = En hårdare variation av ^ trillium ^ där utrymmen endast får fyllas med kungar.
rules.limited.description = Liksom ^ fyrtiofemar ^, men med en 12 av 3 bordau.
rules.lincolngreens.description = En fyrdäcksvariation av ^ puttputt ^ eller en version av ^ panthercreek ^ som tillåter omslagning.
rules.links.description = Ett par-borttagningsspel av Thomas Warfield, avlägset relaterat till ^ golf ^.
rules.linus.description = En lättare variant av ^ labellelucie ^ där du bygger in alternativa färger.
rules.littlebillie.description = I det här spelet som går tillbaka till omkring 1900 är ingen byggnad tillåten, men du har några celler som kan användas för att upptäcka de kort du behöver.
rules.littleforty.description = Liksom ^ fortythieves ^, men vi bygger in oberoende av färg, kan flytta sekvenser och kan göra tre passerar genom däcket och hantera tre kort i taget.
rules.littlegiant.description = En en-däckversion av Giant.
rules.littlemilligan.description = En svåra att vinna en däckversion av ^ missmilligan ^.
rules.littlenapoleon.description = A ^ fortythieves ^ variant som visar några ^ spider ^ influenser, för att du kan bygga oavsett kostym, men bara flytta same-suit sekvenser.
rules.loveaduck.description = A ^ yukon ^ -typ spel, spelat på en sammankopplande bordau.
rules.lower48.description = En variation av ^ fyrtioåtstående ^ där du bygger in alternativa färger istället för i samma färg.
rules.lucas.description = A ^ fortythieves ^ variant med tretton tableau högar och ess som börjar på grunden.
rules.lucasleaps.description = En lätt ^ fortythieves ^ variant som liknar ^ waningmoon ^ förutom att sekvenser kan flyttas.
rules.luckierthirteen.description = En lättare version av ^ luckythirteen ^, eller en cellfri version av ^ freecell ^.
rules.luckyfan.description = En version av ^ freefan ^ där ingen fläkt kan innehålla mer än tre kort.
rules.luckypiles.description = En väldigt lättare variant av ^ Luckythirteen ^ där du kan bygga upp eller ner.
rules.luckythirteen.description = Ett sällan-winnable spel med enkla \
rules.malmaison.description = En svår fyrdäcksversion av ^ josephine ^, eller, om du föredrar, en version av ^ eightythieves ^ som tillåter att sekvenser flyttas.
rules.mamysusan.description = A ^ fortythieves ^ variation från Frankrike med en fem-kort reservera.
rules.manx.description = Bygg färdiga sekvenser genom att omarrangera fyra högar oavsett kostym i detta spel uppfunnet av Rick Holzgrafe of Solitaire Til Dawn.
rules.maria.description = Liksom ^ fyrtiofle ^, men med en 9 till 4 bordau där du bygger i alternerande färger.
rules.marierose.description = En tre-däckversion av ^ josephine ^ eller en version av ^ sexttiotvier ^ som tillåter att sekvenser flyttas.
rules.martha.description = En lätt spel utan lager där halva korten börjar vända neråt.
rules.mcclellan.description = En hårdare variation av ^ littlenapoleon ^ där du behöver bygga i kostym.
rules.midnightclover.description = A ^ fan ^ variant av Thomas Warfield där en rita är tillåten.
rules.midshipman.description = En något lättare variant av ^ maria ^ där vi bygger olika drag i stället för alternativa färger och där några kort börjar utifrån.
rules.millie.description = ^ missmilligan ^ utan reserv.
rules.milligancell.description = A ^ freecell ^ ish variation av ^ missmilligan ^.
rules.milliganharp.description = Ett kors mellan ^ missmilligan ^ och två-deck ^ klondike ^ varianten kallad Harp.
rules.milliganyukon.description = Ett kors mellan ^ milliganharp ^ och ^ yukon ^.
rules.minerva.description = ^ athena ^ med en ^ canfield ^ -stil reserv läggas till.
rules.missmilligan.description = Börja med ett kort i varje kolumn, bygga upp sekvenser med alternativ färg.
rules.mondospider.description = En ganska svår dubbel-storlek åtta kostym ^ spider ^ variant.
rules.moosehide.description = En variant av ^ yukon ^ där du bygger ner i icke-matchande kostymer
rules.morehead.description = A ^ somerset ^ variant där vi bygger olika drag i stället för alternativa färger.
rules.mountolympus.description = Bygg i två år, så odds och evens finns i separata sekvenser på bordet och separata högar på grunden.
rules.movingleft.description = En variant av ^ gargantua ^ eller ^ doubleklondike ^ där tomma utrymmen fylls automatiskt från nästa kolumn.
rules.munger.description = En variation av ^ minerva ^ med reserven är mindre och endast en passerar genom lagret är tillåtet.
rules.muse.description = Denna variation av ^ kingalbert ^ har celler i stället för en reserv.
rules.mystique.description = En variation av ^ munger ^ och ^ minerva ^ med en reserv medelst halvvägs mellan de två.
rules.napoleonsquadrilateral.description = Den här äldre, svårare versionen av ^ napoleonssquare ^ tillåter inte stackförflyttningar, men flyttar mycket kort till grunden under affären.
rules.napoleonsshoulder.description = En varig av ^ napoleonssquare ^ där du bygger oberoende av kostym.
rules.napoleonssquare.description = Detta franska spel, som först beskrivs av Lady Adelaide Cadogen i början av 1900-talet, är en lätt variant av ^ fortythieves ^.
rules.nationale.description = Gilla ^ caprice ^ utan ett lager.
rules.needle.description = Ett spel med en U-formad bordau och en reserv som du kan lagra kort i.
rules.neptune.description = Ett spel där du tar bort par på varandra följande kort.
rules.nestor.description = Kassera några kort med samma rang, oavsett kostym (till exempel två ess, två fiver, etc.).
rules.newyork.description = I den här variationen av ^ dover ^ kan du välja vilken av de tre avfallsspelarna du spelar kort från lageret på, vilket är bra för att det är svårt att omorganisera saker mycket på bordet.
rules.nines.description = En variation på ^ simplepairs ^ par som lägger till 9 eller uppsättning tio genom kung.
rules.northwestterritory.description = Ett kors mellan ^ flowergarden ^ och ^ klondike ^, något lättare än det liknande ^ klondiketerritory ^ spelet.
rules.numberten.description = Liksom ^ fortythieves ^, men två kort i varje tableau-stack hanteras med ansiktet nedåt, vi bygger in alternerande färger och kan flytta staplar som helhet.
rules.octupleklondike.description = En åtta-däck variant av ^ klondike ^.
rules.oddandeven.description = Ett svårt, gammalt och anmärkningsvärt dumt spel där grundstaplar byggs upp i två och ingen byggnad är tillåten på bordet.
rules.odessa.description = En variant av ^ ryska ^ med en annan startbordsbana.
rules.oldcarlton.description = En två-däck ^ klondike ^ -variation, mycket lättare än ^ carlton ^.
rules.opus.description = Thomas Warfields mycket svårare version av ^ pingvin ^ har två färre celler
rules.outback.description = En tvådäcksversion av australiensisk kabal.
rules.pantagruel.description = Denna två-däck ^ klondike ^ -variant är svårare än ^ gargantua ^, men är fortfarande ganska lätt.
rules.panthercreek.description = En fyra-däck ^ golf ^ -variation.
rules.parliament.description = En enklare version av ^ kongressen ^, där esserna börjar på grunden.
rules.passeul.description = A ^ klondike ^ variant med en rektangulär bordau, som skiljer sig från ^ blindalleys ^ endast i antalet passerar genom det tillåtna däcket.
rules.patientpairs.description = Som i ^ simplepairs ^ tar du bort kort med samma rang, men korten börjar utgå till bordet, så en smidgeon är mer skicklig.
rules.penelopesweb.description = En mycket svår variant av ^ beleagueredcastle ^ där utrymmen endast kan fyllas av kungar.
rules.penguin.description = Ett tillfredsställande spel med sju celler som utvecklats av David Parlett, där ett av de kort du behöver för att starta grunden är alltid begravd längst ner i den första bordsskivan.
rules.penta.description = En annan ^ upptagen ^ variation av Thomas Warfield, i den här halvan av tabeau byggs upp och halva bygger ner.
rules.perseverancea.description = En variation av ^ grymt ^ där staplar kan flyttas.
rules.perseveranceb.description = En alternativ version av ^ perseverancea ^ där det bara finns två lösningar, är redningsmetoden annorlunda, och kungar flyttas automatiskt till bottnen av sina staplar.
rules.pharaohs.description = En variation av ^ pyramid ^ med tre pyramider.
rules.phoenix.description = En svårare variant av ^ arizona ^ där du bygger av alternativa färger.
rules.pileup.description = Ett spel där du måste sortera korten genom att rangera istället för att passa.
rules.pitchfork.description = Thomas Warfields variation av ^ nål ^ och ^ höstack ^ där du inte kan bygga på reserven.
rules.pokersquares.description = Gör tio fem-kort pokerhänder från ett 5x5 rutnät.
rules.portuguese.description = En variant av ^ bakersdozen ^ som tillåter att fylla i utrymmen med kungar.
rules.preference.description = En lite mer utmanande version av ^ fortunesfavor ^ med färre tableau högar.
rules.privatelane.description = En variation av ^ beleagueredcastle ^ med två ^ freecell ^ -style-celler tillsattes.
rules.puttputt.description = En lättare variation av ^ golf ^ där inslagning från kung till ess är tillåtet.
rules.pyramid.description = Ett klassiskt parbortspel med en triangulär bordau.
rules.pyramiddozen.description = En version av ^ giza ^ i vilken kort tas bort i par som lägger till tolv.
rules.quadrangle.description = En variation av ^ corona ^ där baskortet bestäms av ett kort som delas in i fundamentet.
rules.quadrennial.description = En version av ^ leapyear ^ med två lösningar eller en version av ^ bekantskap ^ med fyra däck.
rules.quadruplecanfield.description = En enkel fyrdäcksversion av ^ canfield ^ uppfunnad av Thomas Warfield.
rules.quadrupleinterchange.description = En fyrdäcksversion av ^ utbyte ^.
rules.quadrupleklondike.description = En fyrdäcksvariation av ^ klondike ^, uppfunnad av Thomas Warfield.
rules.quadrupletrigon.description = En fyrdäcksversion av ^ trigon ^.
rules.quadrupleyukon.description = En fyrdäcksvariation av ^ yukon ^
rules.queenie.description = Bygga staplar av kort i alternerande färger som i klondike ^, flytta godtyckliga korttyper som i yukon ^ och hantera vågor av kort på bordet, som i ^ spider ^.
rules.queenvictoria.description = Denna mycket lättare variant av ^ kingalbert ^ tillåter att staplar av kort flyttas.
rules.quintupleklondike.description = En fem-däck variant av ^ klondike ^.
rules.quizzie.description = En variation av ^ inquisitor ^ av Thomas Warfield där du hanterar färre kort i varje passera genom däck.
rules.racingaces.description = En tre-deck version av ^ acesandkings ^ uppfunnit av Thomas Warfield.
rules.raglan.description = Detta är ^ kingalbert ^ med en annan tabellau och esser som redan finns på grunden.
rules.rainbow.description = En variation av ^ canfield ^ där du kan bygga oavsett kostym.
rules.rainbowfan.description = Ett dubbelriktat byggnadsspel där du kan rotera kort i staplarna tre gånger.
rules.rankandfile.description = Liksom ^ numren ^, men tre kort i varje stapel behandlas med ansiktet nedåt.
rules.redandblack.description = Ett spel där allt är byggt i alternativa färger.
rules.repair.description = En två-däckversion av ^ freecell ^.
rules.ripplefan.description = En lättare variation av ^ grymt ^ med en ytterligare tabellauhög.
rules.robert.description = Ett nästan oanvändbart spel utan bordläggning.
rules.robie.description = Thomas Warfields version av ^ fortythieves ^ där tableauen börjar tom.
rules.roman.description = En variation av ^ signora ^ där vi bygger oberoende av kostym.
rules.roosevelt.description = En mycket hard ^ fortythieves ^ variant där vi bygger av alternativa färger på bara sju tableau högar.
rules.rougeetnoir.description = En variant av ^ diavolo ^ med en annan tabellau och inget avfall.
rules.rougeforty.description = En variation av ^ rougeetnoir ^ med en rektangulär tabellau.
rules.rowsoffour.description = En enklare version av Diplomat, vilket tillåter vissa lösningar.
rules.royalcotillion.description = En variation av ^ oddandeven ^ med lite extra tableau och reservpiles, men endast ett pass tillåtet genom däck.
rules.royalfamily.description = Det här spelet gör att du kan bygga upp och ner och fylla utrymmen med vilket kort som helst, vilket gör spelet så enkelt att du ofta inte behöver den upplösning som du är tillåten.
rules.royalrendezvous.description = Ett udda österrikiska spel med fyra grundsatser, en normal, en för evens, en för odds och en för kungar.
rules.rueil.description = En version av ^ malmaison ^ underlättades genom att tillåta en redaktion.
rules.russian.description = En hårdare variation av ^ yukon ^ där du måste bygga i samma kostym istället för i alternativa färger.
rules.russiancell.description = Thomas Warfields variant av ^ russian ^ Solitaire lägger till ett par celler.
rules.sally.description = En version av ^ doubleklondike ^ där stiftelsens baskort beror på ett kort som delats in.
rules.sandbox.description = Ett pågående arbete ...
rules.sandboxb.description = Ett annat arbete pågår ...
rules.sanjuanhill.description = En lättare variant av ^ fortythieves ^ där ess redan finns på grunden.
rules.saratoga.description = Det här är bara ^ klondike ^ med korten behandlade med ansiktet uppåt.
rules.sarlacc.description = A ^ freecell ^ variant med en tabellau av interlocking kolumner.
rules.saxony.description = Du har fyra celler, fyra reserverhögar där du kan bygga ner i kostym och åtta bordauhögar, där kort hanteras, men ingen byggnad är tillåten.
rules.scorpion.description = Ett spel med en sju-i-sju bordau, där tre kort i de fyra första staplarna börjar vända neråt.
rules.scorpionhead.description = En variation av ^ scorpion ^ med några celler.
rules.scorpiontail.description = En variant av ^ scorpion ^ där vi bygger ner med alternativ färg i stället för ner i kostym.
rules.scotch.description = Stiftelser bygger i alternativa färger, bordau bygger oavsett kostym.
rules.seatowers.description = En populär ^ freecell ^ -variation uppfunnad 1988 av Art Cabral.
rules.selectivecastle.description = En version av ^ beleagueredcastle ^ där basen av grunden bestäms av det första kortet du spelar för det.
rules.selectivefreecell.description = En variation av ^ freecell ^ där det första kortet spelade till foudnation sätter grundvärdet för alla fundamenten.
rules.sevastopol.description = En enklare version av ^ kiev ^ där fyra bordauhögar börjar med tre kort istället för fyra.
rules.sevenbyfive.description = A ^ freecell ^ variant med en mindre tabellau kolonn och mer mer cell.
rules.sevenbyfour.description = En hårdare ^ freecell ^ variant med en mindre tabellau kolonn.
rules.sevenbyseven.description = Detta danska spel med en sju-i-sju tabellau och tre celler tillåter två redes.
rules.sevendevils.description = Sju Devils är förmodligen det svåraste av alla solitaire-spel.
rules.sextupleklondike.description = En sex-däck variant av ^ klondike ^.
rules.shadylanes.description = Ett svårt spel med fyra reserverhögar och fyra bordauhögar.
rules.shamrocks.description = En variation av ^ fan ^ där du kan bygga upp eller ner oberoende av kostym, men är begränsade till tre kort per stapel.
rules.shuffle.description = En version av ^ neptune ^ där du också kan para konungar med ess.
rules.signora.description = Bygg allt i alternativa färger, samtidigt som du försöker rensa en elva kort reserv till Foundaton.
rules.simonjester.description = En två-däck variant av ^ simplesimon ^ uppfunnad av Adam Selene.
rules.simonsays.description = En blandning av ^ simplesimon ^ med ^ freecell ^ uppfunnad av Thomas Warfield.
rules.simplepairs.description = Ett spel där du tar bort kort med samma rang.
rules.simplesimon.description = Liksom en däck ^ spindel ^ där alla kort börjar vända upp i en triangulär bordau och det finns inga ytterligare kort att hantera.
rules.singleinterchange.description = En svår en-däckvariant av ^ utbyte ^ uppfunnet av Thomas Warfield.
rules.singleleft.description = Thomas Warfields en-däckversion av ^ movingleft ^.
rules.singlerail.description = En däckversion av ^ doublerail ^.
rules.sirtommy.description = Ett klassiskt gammalt solitaire spel där kort kan placeras var som helst på bordet, men kan inte omorganiseras.
rules.sixbyfour.description = En mycket hårdare ^ freecell ^ variant med två färre tabellau kolumner.
rules.sixesandsevens.description = Ingen byggnad på bordau, någon grundbyggnad byggs upp, vissa bygger sig ner.
rules.sixteenpiles.description = Ett ovanligt spel där du staplar kort med samma nivåer för att ta fram kort för att flytta till grunden.
rules.sixtythieves.description = En svår tre-deck version av ^ fortythieves ^ av Thomas Warfield.
rules.skippy.description = Ett spel uppfunnet av Lillian Davies och Christa Baran.
rules.smokey.description = A ^ klondike ^ variant uppfunnad av Ann Edwards där du kan bygga sekvenser i färg, men bara flytta sekvenser av samma färg.
rules.somerset.description = A ^ klondike ^ variant utan lager eller avfall.
rules.spanish.description = En variant av ^ bakersdozen ^ som tillåter att fylla i utrymmen.
rules.spider.description = På de 10 bordau-staplarna kan du bygga ner oavsett kostym, men du kan bara flytta enkla kostsekvenser.
rules.spidercells.description = A ^ freecell ^ variant där du behöver bygga fullständiga växlande färgsekvenser på bordet.
rules.spiderette.description = En en-däckversion av ^ spider ^, med en ^ klondike ^ -stil triangulär tabellau.
rules.spideronesuit.description = ^ Spider ^ med ingenting annat än spader, spader, spader, så långt ögat kan se.
rules.spiderthreedeck.description = Denna tre-däckversion av ^ spider ^ är lite lättare än ^ bigspider ^.
rules.spidertwosuits.description = Namnet säger det \
rules.spidike.description = Thomas Warfields blandning av ^ spider ^ med en ^ klondike ^ slutar ser mycket ut som ^ spiderette ^ förutom att kort kan flyttas enstaka till grunden.
rules.spike.description = ^ klondike ^ med tre avfallspiller.
rules.squadron.description = En mycket lättare version av ^ fortythieves ^ med tre celler.
rules.stages.description = En lättare variant av ^ upptagssatser ^ som tillåter stapelrörelser.
rules.stalactites.description = Det här otroliga spelet utan byggnad kräver att du rensar bordau med bara två celler som hjälper dig.
rules.steps.description = En två-däckversion av ^ klondike ^.
rules.steve.description = En två-däck ^ klondike ^ variant där vi bygger oberoende av kostym, men kan bara flytta samma kostymsekvenser.
rules.stewart.description = En svårare variation av ^ martha ^ i vilken endast enstaka kort kan flyttas.
rules.stonewall.description = På samma sätt som ^ flowergarden ^, förutom att vissa kort börjar vända ner, måste du bygga in alternativa färger, och du kan flytta sekvenser.
rules.storehouse.description = En gammal ^ canfield ^ -variant som först beskrivits 1939. Ett trevligt spel, men det behövs knappast någon strategi.
rules.straightfifteens.description = En lättare variation av ^ fiftefen ^ där tiotals, jacks, queens och kungar avlägsnas i grupper som innehåller en av varje i stället för fyra i ett slag.
rules.strata.description = En åtta-åtta kvadratisk bordau, en kort däck och två lösningar gör det här spelet intressant.
rules.streets.description = Precis som ^ fortythieves ^, förutom att du bygger in alternativa färger.
rules.streetsandalleys.description = En svårare variation av ^ beleagueredcastle ^ som börjar med inga kort som delas in i stiftelsen.
rules.stronghold.description = En variant av ^ beleagueredcastle ^ med en ^ ^ freecell ^ stilcell tillsattes.
rules.suitelevens.description = En variation av ^ elevens ^ där du bara kan ta bort uppsättningar kort om de är alla av samma färg.
rules.suitsup.description = En enkel match där du tar bort kort av samma färg, tills endast fyra kort är kvar.
rules.suittriangle.description = En två-däckversion av ^ klondike ^ där vi bygger i samma svit.
rules.superchallengefreecell.description = En version av ^ freecell ^ uppfunnad av Thomas Warfield där ess och twos alltid ligger på botten av de åtta staplarna och där utrymmen endast kan fyllas av kungar.
rules.superflowergarden.description = Det här är en enklare version av ^ märkellucus ^ i vilken man kan bygga oavsett kostym.
rules.superiorcanfield.description = Canfield gjorde lite lättare och lite mer strategiskt genom att hantera reservkorten och vända sig inte automatiskt till reserven.
rules.sweetsixteen.description = En variant av ^ trustytwelve ^ där du bygger av alternativ färg
rules.swiss.description = Liksom ^ klondike ^ men essar är höga och tableauen är pyramidisk.
rules.tabbycat.description = En enklare version av ^ manx ^ som tillåter en sekvens att parkeras i svansen.
rules.takingsilk.description = En två däckversion av ^ thirtysix ^.
rules.tarantula.description = En lättare variant av ^ spider ^ där du får flytta sekvenser som alla är en färg även om de inte är alla ena kostym.
rules.tenacross.description = En variation av ^ ryska ^ med en annan start tabell och två celler, som börjar vara fulla.
rules.tenbyone.description = Tio tableau-staplar och en cell gör ett spel med likheter med ^ freecell ^ och ^ vingård ^.
rules.tens.description = Ett uppsättning avlägsningsspel som liknar ^ simplepairs ^ där du kan ta av par som lägger till 10 eller en uppsättning fyra matchande kort tio eller högre.
rules.tensout.description = En variation av ^ fourteenout ^ där vi tar bort par som lägger till 10.
rules.thewish.description = Detta enkla parborttagningsspel använder en kort däck och inget lager, men liknar annars ^ dubblets ^.
rules.thievesofegypt.description = En variant av ^ fortythieves ^ med en pyramidformad tableau.
rules.thievesrush.description = A ^ fortythieves ^ variant uppfann av Thomas Warfield där i var och en passerar genom däcken du hanterar i mindre bitar.
rules.thirteens.description = Ta bort par som lägger till tretten.
rules.thirtyninesteps.description = ^ waningmoon ^ med färre kort i den ursprungliga tabellen.
rules.thirtysix.description = En sex-i-sex tabellau där du bygger oberoende av färg.
rules.thoughtful.description = ^ klondike ^ med alla kort i bordet börjar uppifrån.
rules.threebears.description = En variation på ^ tripleklondike ^ uppfunnad av Thomas Warfield.
rules.threeblindmice.description = En variation av ^ scorpion ^ med en 10 till 5 bordau och en två-kort reserv.
rules.threecell.description = En variation av ^ freecell ^ med endast tre celler.
rules.threedemons.description = Denna tre-däckversion av ^ canfield ^ som uppfunnits av Thomas Warfield börjar med flera kort i reserven och fler bordauhögar än ^ triplecanfield ^.
rules.threepirates.description = En variation av ^ fyrtiofle ^ med tre avfallspiller.
rules.threescompany.description = En ganska svår variant av ^ deuces ^ eller ^ busyaces ^ med ännu färre tableau högar men stack flyttningar är tillåtna.
rules.threeshufflesandadraw.description = En variation av ^ märkljus ^ som lägger till en rita.
rules.thumbandpouch.description = Liksom ^ klondike ^, men lättare, eftersom kort kan spelas på bordau kort av någon annan kostym.
rules.titan.description = En version av ^ jätte ^ som börjar med fler kort på bordet.
rules.tournament.description = Ett tvådäcksspel där ingen byggnad är tillåten på bordet, och du måste förlita dig åt åtta celler för att flytta dina kort till grunden.
rules.trefoil.description = En något lättare variation av ^ märkellucus ^ där esserna börjar på grunden och det finns färre tabellau kolumner.
rules.trevigarden.description = En variation av ^ stonewall ^ underlättades genom tillsats av två celler.
rules.triangle.description = En mycket svår inverterad version av ^ pyramid ^.
rules.trigon.description = En variation av ^ klondike ^ där vi bygger in kostym istället för med växlande färger.
rules.trigonleft.description = En blandning av ^ trigon ^ och ^ movingleft ^.
rules.trillium.description = A ^ spider ^ variant med en 13x4 bordau där du bygger ner efter alternativ färg.
rules.triplecanfield.description = En lätt tre-däckversion av ^ canfield ^ uppfunnad av Thomas Warfield som har färre bordshögar och en mindre reserv än ^ treemder ^.
rules.tripleeasthaven.description = En tre-däckversion av ^ easthaven ^ av Thomas Warfield.
rules.triplefourteens.description = En tre-däckversion av ^ fourteenout ^ som uppfanns av Thomas Warfield.
rules.triplefreecell.description = Thomas Warfields tre-däckversion av ^ freecell ^.
rules.tripleharp.description = En tre-däckversion av ^ harp ^ uppfunnad av Thomas Warfield.
rules.tripleinterchange.description = En tre-däckversion av ^ utbyte ^.
rules.tripleklondike.description = En tre däckversion av ^ klondike ^ uppfunnad av Thomas Warfield.
rules.tripleleft.description = Thomas Warfields tre-däckversion av ^ movingleft ^.
rules.tripleminerva.description = Thomas Warfields tre-däckversion av ^ minerva ^.
rules.triplerussian.description = En tre-däckversion av ^ russian ^ solitaire av Thomas Warfield.
rules.triplescorpion.description = En tre-däck variant av ^ scorpion ^ utan reserv.
rules.tripletriangle.description = En tre-deck ^ eternaltriangle ^ variation av Thomas Warfield.
rules.tripleyukon.description = En tre-däckvariation av ^ yukon ^
rules.trustytwelve.description = Mer lycka än färdighet behövs för att vinna detta spel byggsekvenser på bordet.
rules.tuxedo.description = En lättare variant av ^ pingvin ^ där alla kort börjar på bordet.
rules.tvetesgrandfather.description = Paul Olav Tvete lärde sig detta spel från sin farfar och inkluderade det i KPatience.
rules.twenty.description = Ett något meningslöst spel med tjugo reserverhögar och ingen byggnad.
rules.twocell.description = En variation av ^ freecell ^ med endast två celler.
rules.ukrainian.description = En sällan winnable version av ^ russian ^ Solitaire där endast fullständiga sekvenser kan tas bort, som i spindel.
rules.unlimited.description = En lättare variant av ^ utbyte ^, där vi får obegränsade förklaringar
rules.unusual.description = En två-däckversion av ^ grym ^.
rules.upandup.description = En variation av ^ trustytwelve ^ där du kan bygga kungar på ess.
rules.usk.description = A ^ klondike ^ variant utan lager eller avfall.
rules.variegatedcanfield.description = En svår tvådäcksversion av ^ canfield ^, med ess som börjar på grunden och endast tre passerar genom det tillåtna avfallet.
rules.vineyard.description = En svår variant av ^ bakersdozen ^ uppfunnad av Peter Voke.
rules.wadingpool.description = En lättare variation av ^ wavemotion ^ som tillåter att bygga, men inte stapla rörelser, på reserven.
rules.waningmoon.description = A ^ fortythieves ^ variant med fler tableau högar.
rules.waterloo.description = A ^ fortythieves ^ variant med ^ spider ^ -liknande byggregler.
rules.wavemotion.description = I David Bernazzani''s variation på ^ freecell ^ och ^ scorpion ^ börjar alla kort på reserven.
rules.waxingmoon.description = En mycket svår ^ förtythieves ^ variant av Thomas Warfield.
rules.westcliff.description = En väldigt lätt ^ klondike ^ variant där du har tio tableau högar.
rules.whitehead.description = Liksom ^ klondike ^, men med kort vänd uppåt och du bygger i matchande färger i stället för alternerande färger.
rules.whitehorse.description = En enkel ^ klondike ^ variant där vi istället för att hantera mycket kort till bordet har utrymmen som autofyller
rules.wildflower.description = En variation av ^ flowergarden ^ där du kan flytta sekvenser av kort i samma färg tillsammans.
rules.willothewisp.description = En däckversion av ^ spider ^, med en rektangulär 7x3 bordau.
rules.willow.description = A ^ klondike ^ -variation med fyra fanhögar där vi kan bygga med kort med samma rang.
rules.winery.description = En version av ^ vingård ^ med celler tillsattes.
rules.wood.description = Ett spel där vi bygger både grunden och bordet i alternativa färger.
rules.yakutatbay.description = Ett kors mellan ^ yukon ^ och ^ movingleft ^.
rules.yukon.description = Ett välkänt spel med inget lager, där staplar av kort kan flyttas även om de inte är i följd.
rules.yukoncells.description = En variation av ^ yukon ^ förenklas genom tillsatsen av två celler.
rules.yukonicplague.description = En svårare variation av ^ yukon ^ där många kort är begravda i en reserv.
rules.yukonkings.description = En svår version av ^ yukon ^ utan stiftelser.
rules.yukononesuit.description = En en-kostvariation av ^ yukon ^.
rules.zerline.description = Ett tyskt spel där drottningar är höga och du har en kortplats för fyra kort.